module main();
    // Typewriter mechanical logic
    typewriter tw();
endmodule
